package shared_pkg;
    parameter WRITE_LOOP = 5;
    parameter READ_LOOP = 5;
endpackage